module mux16(input wire [0:15] i, input wire [3:0] j, output wire o);
	wire  t0, t1;
	mux8 mux8_0 (i[0:7], j[0], j[1], j[2], t0);
	mux8 mux8_1 (i[8:15], j[0], j[1], j[2], t1);
	mux2 mux2_0 (t0, t1, j[3], o);
endmodule

module left_shift(input wire [15:0] i, input wire [3:0] shift, output wire [15:0] o);
	mux16 mux16_15( { i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0] }, shift, o[15]);
    mux16 mux16_14( { i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0 }, shift, o[14]);
    mux16 mux16_13( { i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0 }, shift, o[13]);
    mux16 mux16_12( { i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0 }, shift, o[12]);
    mux16 mux16_11( { i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[11]);
    mux16 mux16_10( { i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[10]);
    mux16 mux16_9( { i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[9]);
    mux16 mux16_8( { i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[8]);
    mux16 mux16_7( { i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[7]);
    mux16 mux16_6( { i[6], i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[6]);
    mux16 mux16_5( { i[5], i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[5]);
    mux16 mux16_4( { i[4], i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[4]);
    mux16 mux16_3( { i[3], i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[3]);
    mux16 mux16_2( { i[2], i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[2]);
    mux16 mux16_1( { i[1], i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[1]);
    mux16 mux16_0( { i[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[0]);
endmodule

module right_shift(input wire [15:0] i, input wire [3:0] shift, output wire [15:0] o);
	mux16 mux16_0( { i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15] }, shift, o[0]);
    mux16 mux16_1( { i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0 }, shift, o[1]);
    mux16 mux16_2( { i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0 }, shift, o[2]);
    mux16 mux16_3( { i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0 }, shift, o[3]);
    mux16 mux16_4( { i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[4]);
    mux16 mux16_5( { i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[5]);
    mux16 mux16_6( { i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[6]);
    mux16 mux16_7( { i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[7]);
    mux16 mux16_8( { i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[8]);
    mux16 mux16_9( { i[9], i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[9]);
    mux16 mux16_10( { i[10], i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[10]);
    mux16 mux16_11( { i[11], i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[11]);
    mux16 mux16_12( { i[12], i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[12]);
    mux16 mux16_13( { i[13], i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[13]);
    mux16 mux16_14( { i[14], i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[14]);
    mux16 mux16_15( { i[15], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }, shift, o[15]);
endmodule

module left_rotate(input wire [15:0] i, input wire [3:0] shift, output wire [15:0] o);
	mux16 mux16_15( { i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0] }, shift, o[15]);
    mux16 mux16_14( { i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15]}, shift, o[14]);
    mux16 mux16_13( { i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14] }, shift, o[13]);
    mux16 mux16_12( { i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13] }, shift, o[12]);
    mux16 mux16_11( { i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12] }, shift, o[11]);
    mux16 mux16_10( { i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11] }, shift, o[10]);
    mux16 mux16_9( { i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10] }, shift, o[9]);
    mux16 mux16_8( { i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9] }, shift, o[8]);
    mux16 mux16_7( { i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8] }, shift, o[7]);
    mux16 mux16_6( { i[6], i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7] }, shift, o[6]);
    mux16 mux16_5( { i[5], i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6] }, shift, o[5]);
    mux16 mux16_4( { i[4], i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5] }, shift, o[4]);
    mux16 mux16_3( { i[3], i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4] }, shift, o[3]);
    mux16 mux16_2( { i[2], i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3] }, shift, o[2]);
    mux16 mux16_1( { i[1], i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2] }, shift, o[1]);
    mux16 mux16_0( { i[0], i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1] }, shift, o[0]);
endmodule

module right_rotate(input wire [15:0] i, input wire [3:0] shift, output wire [15:0] o);
	mux16 mux16_0( { i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15] }, shift, o[0]);
    mux16 mux16_1( { i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0] }, shift, o[1]);
    mux16 mux16_2( { i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1] }, shift, o[2]);
    mux16 mux16_3( { i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2] }, shift, o[3]);
    mux16 mux16_4( { i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3] }, shift, o[4]);
    mux16 mux16_5( { i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4] }, shift, o[5]);
    mux16 mux16_6( { i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5] }, shift, o[6]);
    mux16 mux16_7( { i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6] }, shift, o[7]);
    mux16 mux16_8( { i[8], i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7] }, shift, o[8]);
    mux16 mux16_9( { i[9], i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8] }, shift, o[9]);
    mux16 mux16_10( { i[10], i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8],i[9] }, shift, o[10]);
    mux16 mux16_11( { i[11], i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10] }, shift, o[11]);
    mux16 mux16_12( { i[12], i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11] }, shift, o[12]);
    mux16 mux16_13( { i[13], i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12] }, shift, o[13]);
    mux16 mux16_14( { i[14], i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13] }, shift, o[14]);
    mux16 mux16_15( { i[15], i[0], i[1], i[2], i[3], i[4], i[5], i[6], i[7], i[8], i[9], i[10], i[11], i[12], i[13], i[14] }, shift, o[15]);
endmodule

module alu(input wire [15:0] i, input wire [3:0] shift, input wire [1:0] op, output wire [15:0] o);
	wire [15:0] o_ls, o_rs, o_lr, o_rr;
	left_shift ls_0(i, shift, o_ls);
	right_shift rs_0(i, shift, o_rs);
	left_rotate lr_0(i, shift, o_lr);
	right_rotate rr_0(i, shift, o_rr);

	assign o = (op[1] == 1'b0) ? ((op[0] == 1'b0) ? o_ls : o_rs) : ((op[0] == 1'b0) ? o_lr : o_rr);

endmodule